`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:21:32 06/15/2022 
// Design Name: 
// Module Name:    InstructionMemory 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module InstructionMemory(
		address, inst
    );
	
	input [19:0] address;
	output reg [19:0] inst;
		
	reg [19:0] mem [31:0];
	
	always @ (*)
	begin
	mem[0] = 20'b00000000000000000000;  
   mem[1] = 20'b00000000000000000001;  
   mem[2] = 20'b00000000000000000010;  
   mem[3] = 20'b00000000000000000011;  
   mem[4] = 20'b00000000000000000100;  
   mem[5] = 20'b00000000000000000101; 
   mem[6] = 20'b00000000000000000110;  
   mem[7] = 20'b00000000000000000111;  
	
   mem[8] = 20'b00000000000000000000;  
   mem[9] = 20'b00000000000000000000;  
   mem[10] = 20'b00000000000000000000;  
   mem[11] = 20'b00000000000000000000;  
   mem[12] = 20'b00000000000000000000;  
   mem[13] = 20'b00000000000000000000;  
   mem[14] = 20'b00000000000000000000;  
   mem[15] = 20'b00000000000000000000;
	
 	mem[16] = 20'b00001000000110000000;  
   mem[17] = 20'b00000010110010110010;  
   mem[18] = 20'b00001101110001100111;  
   mem[19] = 20'b00001101110111011001;  
   mem[20] = 20'b00001111110110110001;  
   mem[21] = 20'b00001100000001111011; 
   mem[22] = 20'b00000000000000000000;  
   mem[23] = 20'b00000000000000000000;
	
   mem[24] = 20'b00000000000000000000;  
   mem[25] = 20'b00000000000000000000;  
   mem[26] = 20'b00000000000000000000;  
   mem[27] = 20'b00000000000000000000;  
   mem[28] = 20'b00000000000000000000;  
   mem[29] = 20'b00000000000000000000;  
   mem[30] = 20'b00000000000000000000;  
   mem[31] = 20'b00000000000000000000; 
	
	inst = mem[address[4:0]];
	end
	
	

endmodule
